library verilog;
use verilog.vl_types.all;
entity al422b_2rgb_8s_vlg_tst is
end al422b_2rgb_8s_vlg_tst;
